// Code your design here
module encoder(s,y);
  input[3:0]s;
  output reg [1:0]y;
  always@(*)begin
    case(s)
      4'b0001:y=2'b00;
      4'b0010:y=2'b01;
      4'b0100:y=2'b10;
      4'b1000:y=2'b11;
      default:y=2'b00;
    endcase
  end
endmodule

interface inter;
  logic[3:0] s;
  logic[1:0] y;
endinterface
