//constraint == means restruction
//solve before constraint:
class sample;
  rand bit[7:0]a,b;
  constraint c1{solve a before b;}
  constraint c2{ b==a-15;}
endclass

module tb;
  sample s=new();
  initial begin
    assert(s.randomize());
    $display("a=%0d,b=%0d",s.a,s.b);
  end
endmodule
//output:
# KERNEL: a=39,b=24
