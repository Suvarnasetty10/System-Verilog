//Descending order of the array
class sample;
  int i,j;
  rand bit[3:0] a[];
  int val;
  constraint c1 {a.size==10; //element count
                 foreach(a[i]){
                   if(i>0)
                     a[i]<a[i-1];
                }
                }
endclass
module tb;
  sample s=new();
  int i;
  initial begin
    assert(s.randomize());
    foreach(s.a[i])
    $display("a[%0d]=%0d ",i,s.a[i]);   
  end
endmodule
//output:
# KERNEL: a[0]=14 
# KERNEL: a[1]=13 
# KERNEL: a[2]=11 
# KERNEL: a[3]=9 
# KERNEL: a[4]=8 
# KERNEL: a[5]=5 
# KERNEL: a[6]=4 
# KERNEL: a[7]=2 
# KERNEL: a[8]=1 
# KERNEL: a[9]=0 
                 
                 
                 
                 
