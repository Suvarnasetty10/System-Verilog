class parent;
   int a=10;
   int b=7;
  function void print();
    $display(" a=%0d, b=%0d",a,b);
  endfunction
endclass

class child extends parent;
  int c;
  function void sub();
    c=a-b;
    $display(" c=%0d",c);
  endfunction
endclass
 
module tb;
  int d;
  child c;
  initial begin
    c=new();
    c.print();
    c.sub();
  end
endmodule
//output:
# KERNEL:  a=10, b=7
# KERNEL:  c=3




  
  
